library ieee;

entity actividad1 is
    port (
        
    );
end entity actividad1;

architecture rtl of actividad1 is
    
begin
    
    
    
end architecture rtl;